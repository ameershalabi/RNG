--------------------------------------------------------------------------------
-- Title       : casr test vectors inputs/outputs
-- Project     : hdl_rand
--------------------------------------------------------------------------------
-- File        : casr_test_vectors_pkg.vhd
-- Author      : Ameer Shalabi <ameershalabi94@gmail.com>
-- Last update : Fri Jan 16 14:54:05 2026
--------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- Description: casr package with test vectors
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

package casr_test_vectors_pkg is

    constant casr30_seed1_c     : std_logic_vector(63 downto 0)  := x"36BD0F75A4ABE07D";
    constant casr90_seed1_c     : std_logic_vector(127 downto 0) := x"DB33FA5E3C4D8A2C36BD0F75A4ABE07D";
    constant casr150_seed1_c    : std_logic_vector(255 downto 0) := x"FC7FFDD5E74EF4C24F7F1722EF758AC4DB33FA5E3C4D8A2C36BD0F75A4ABE07D";
    constant casr90150h_seed1_c : std_logic_vector(511 downto 0) := x"285F44AB321ED5E5D7F04BB5AD4D5B981EC6F4E08D475D5F8E7DBBB955F6389DFC7FFDD5E74EF4C24F7F1722EF758AC4DB33FA5E3C4D8A2C36BD0F75A4ABE07D";
    constant casr90150h_rule1_c : std_logic_vector(511 downto 0) := x"FC7FFDD5E74EF4C24F7F1722EF758AC4DB33FA5E3C4D8A2C36BD0F75A4ABE07D285F44AB321ED5E5D7F04BB5AD4D5B981EC6F4E08D475D5F8E7DBBB955F6389D";

    constant n_gen_rand : integer := 100;
    type casr30_vectors_t is array (0 to n_gen_rand-1) of std_logic_vector(63 downto 0);
    constant casr30_vectors : casr30_vectors_t := (
            x"D2859114BFA83085",x"5ECCFBB780AC59CC",x"C2770890C1A6CE76",x"67919DF962BA7392",x"B8FAE40F368B9CFF",
            x"8D0A3E11D2D8E700",x"D59B433A5E4D3981",x"54E965CBC3F5CEC2",x"D72F3C7864147267",x"51E1C68CBE369FB8",
            x"DA326AD78352E08C",x"4B5FAA50C55E31D7",x"7940ABD96D435A51",x"0F61A84F25654BDB",x"9132ACF1FD3D7849",
            x"FBDEA71A05C50CFE",x"0842B9AB0C6D9702",x"1CE68EA996A4F187",x"A73AD2AEF2BF1AC9",x"B9CA5EA21E81AA7E",
            x"8E7BC2B722C2AB82",x"D3886691F666A8C6",x"5CDCBAFA13BAAD6A",x"C7478A0B3C8AA52B",x"6968DB19C7DABDE8",
            x"AF2D49AE684A842C",x"A1E57EA3ACFACE67",x"B23D02B4A70A73B8",x"9F458697B99B9C8D",x"E16CCAF08EE8E7D4",
            x"33277A19D22D3857",x"DDF90B2E5F65CCD1",x"440F99E3C13C775A",x"EE10EE3463C6914B",x"23392356B46AFB78",
            x"75CFF55296AA090C",x"9470155EF2AB1F96",x"F69835421EA9A0F2",x"12EC556722AEB11E",x"3E26D539F6A29BA3",
            x"C37A55CE12B6E8B5",x"650BD4733E922D94",x"BD98569DC2FF64F6",x"84ECD2E466013F12",x"CF275E3EBB03C1BE",
            x"71F9434289846282",x"9A0F6566DECEB6C7",x"EB113D3A42729268",x"29BBC5CBE79EFFAD",x"EE886C7838E200A5",
            x"22DCA68C4D3701BC",x"7647BAD6F5D18286",x"93E88A52145AC6CB",x"FC2DDBDF36CA6A78",x"06644841D27BAB8D",
            x"8BBEFCE25F88A8D5",x"D8820737C0DDAD54",x"4DC709D06144A557",x"74699E58B36FBD51",x"16AEE3CD9D20855B",
            x"B2A23474E5F1CD49",x"9EB756973C1A757E",x"E29152F1C62B9502",x"36FB5E1A6B68F586",x"5209432BA92D14CB",
            x"5F1F65E8AFE5B779",x"41A13C2DA03C910F",x"62B3C664B047FB91",x"369C6BBF98E808FB",x"D2E6A880ED2C1D09",
            x"5E3AADC125E6259E",x"C34AA463FC3B7CE3",x"657ABEB406490734",x"BD0A82960BFF89D6",x"859AC6F31800DE52",
            x"CCEA6A1DAC0143DE",x"772BAB24A6036442",x"91E8A9FFBB053EE7",x"FA2DAE00898DC238",x"0B64A301DED4674D",
            x"993FB5824256B975",x"EFC094C7E7D28F14",x"2061F768385ED1B7",x"F0B2112C4CC25A91",x"199F3BE6F767CAFA",
            x"2EE1C83A11387A0B",x"E2327C4B3BCC8B19",x"375F86F9C877D9AE",x"5140CA0E7C904EA3",x"5B617B1387F8F2B5",
            x"493309BCC80D1E95",x"7FDD9E877C15A2F5",x"0044E2C90634B615",x"80EF367F8B579335",x"C121D380D950FDD4",
            x"63F25CC14F590457",x"341FC763714F8ED1",x"D62069351B70D25B",x"5370AFD5A9195FC8",x"DD19A054AFAF407C"
        );

    type casr90_vectors_t is array (0 to n_gen_rand-1) of std_logic_vector(127 downto 0);
    constant casr90_vectors : casr90_vectors_t := (
            x"5BFE099366BDD14E762499519B0230C5",x"1A0317EF7E254A3BD75B7E0BFB8579E8",x"3907A4294358316A451B43120AC84F24",
            x"6E8C9A46271C7A61A8BB27AD10F4B9DA",x"EA5F79AF5DB6C9F3852BDC8CA9932F59",x"21914F8915B6F71EC8C2575F07EFC91F",
            x"D3EA38D6A1B695B2F5E585118C2876B1",x"4E216DC613B661BC9139C8ABDE44D63B",x"3B526D6F2EB7F3A76AEF750253ABC76B",
            x"EB0DEC69CA341E9D60A950858E826D63",x"239D2EE77172327471060949DA45EC76",x"56F4CABD5A5D7DD2DA8F163759A92ED7",
            x"0693F0241994454CD859A7751F86CAC5",x"8E6E185A3FE2A83FDC9F9D50B0CEF0E8",x"5BEB3C99603404605770F40939FA99A5",
            x"1A23E77E70720AF085599216EF087F98",x"39563D43D8DD1099481FED26A994C0FC",x"6E0764265DD4A97E34302CDE07E3E186",
            x"EB0D7A5F9543064372784FD30C3633CF",x"239C4990E0278FA75DCCB84F9E777E78",x"56F6B7E9B05CD89D157F2CB8F3D543CC",
            x"86963427B897DD74A041CF2D9E40267E",x"4E67725CAD64545310A379CDF3A05FC2",x"BBFD5D970C7A828FA9174F7D1E909065",
            x"AA0415E59EC8445886A53944B26968F9",x"810A2139F2F4AA9D4E18EE2B3DE6658F",x"C29152EF1C9300743B3DAB43E53FF9D8",
            x"E46A0CA9B76F80D26BE5832638E00F5D",x"3AE11F07B568C1CDE239C7DF6DB01915",x"E8B2B18CB065E37D356F6C516DB83EA0",
            x"A53C3BDF38F93744F0696E8A6DAC6211",x"98E66A51ED8EF52B98E66A51ED8EF52B",x"FDBFE18B2DDA90C2FDBFE18B2DDA90C2",
            x"85A033D3CD5869E485A033D3CD5869E4",x"49907E4E7C1CE73B49907E4E7C1CE73B",x"37E8C3BBC637BDEB37E8C3BBC637BDEB",
            x"F425E6AA6F74A523F425E6AA6F74A523",x"12593E01E95318D612593E01E95318D6",x"2D9EE303260FBDC72D9EE303260FBDC7",
            x"CDF2B787DF18A56DCDF2B787DF18A56D",x"7D1C34CC51BD186D7D1C34CC51BD186D",x"44B673FE8BA4BCEC44B673FE8BA4BCEC",
            x"AB37DE02529B27AEAB37DE02529B27AE",x"03F453058C7BDC8A03F453058C7BDC8A",x"06128F89DECA575106128F89DECA5751",
            x"8F2C58D752F1850A8F2C58D752F1850A",x"59CE9DC50C9BC89059CE9DC50C9BC890",x"9F7A75689F7A75689F7A75689F7A7568",
            x"7149D0657149D0657149D0657149D065",x"5A3748F85A3748F85A3748F85A3748F8",x"9975358C9975358C9975358C9975358C",
            x"7E50F1DF7E50F1DF7E50F1DF7E50F1DF",x"43899B5143899B5143899B5143899B51",x"26D7FB0A26D7FB0A26D7FB0A26D7FB0A",
            x"5EC40B915EC40B915EC40B915EC40B91",x"12EA12EA12EA12EA12EA12EA12EA12EA",x"2CA12CA12CA12CA12CA12CA12CA12CA1",
            x"CF12CF12CF12CF12CF12CF12CF12CF12",x"F9ACF9ACF9ACF9ACF9ACF9ACF9ACF9AC",x"8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F8F",
            x"D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8D8",x"DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD",x"55555555555555555555555555555555",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000",x"00000000000000000000000000000000",x"00000000000000000000000000000000",
            x"00000000000000000000000000000000"
        );


    type casr150_vectors_t is array (0 to n_gen_rand-1) of std_logic_vector(255 downto 0);
    constant casr150_vectors : casr150_vectors_t := (
            x"FABFF894DA746727F63EB2F646245A2F00CDF3CD5AF05B62409996243FA9D0B8",
            x"729FF5F703A69AFBE15C8E61E97EC3668130EDB14268C017E1E6717E5F2E9995",
            x"2EEFE4E28538E271D34BD592CF3C2418C3C9400B678D2033D2D9AB3DCEE4E675",
            x"E447DF56CDD557AA9C79947E36DA7E2525BF60181B51F04D9E0628D8B45F59A5",
            x"DEEB8E503095532AEAB676BD4003BD7DFC1E1024205AE8F06D096D0586CE463C",
            x"0C4955D849F55CEA4A81A09960051938FA2D387E70C24D68819F018C4835E95B",
            x"92FF5484FEE54B4BFAC231E7100DA7D57361D4BDA927F10DC26E8252FC44CF40",
            x"FE7E57CF7C5D7879F2274ADAB8103B952C1297982FFBEB90A784C7DE7AEF3661",
            x"FDBDD3B63AC934B6EF7A7A0294385175E23EF36467F1C979BB4F2B8DB246C192",
            x"78189D01523FC7804633B306F654DB24D75C6C1E9BEABF361076E9500FE8227E",
            x"B425E9835F5FAB40E94D0C8861D700FF124A822CE1CA9EC138A04F5817CC77BD",
            x"067CCE444E4F28614F7193DC9292817EBFFAC76352BAEC23D5B0F64433B2A318",
            x"09BB35EEF5F6EC93762A7D8BFEFEC33C9FF22A145E924275940961EE4D0EB4A4",
            x"1E10C4C464E043FC216BB859FC7C24DBEFEF6B36CCFFE7A4761F12C5F19487BE",
            x"2D392F2E9F50E5FA730914C6FABA7F01C7C608C0337FDB3EA12EBE2CEA77CB1D",
            x"E1D7E6E4EE595CF3AC9FB7287293BE82ABA91D204C3F80DCB3E49D634BA3B8A9",
            x"D293D85F45C74B6D23EF02ECAEFD1CC6A92FA9F0F25F410B8DDFE914793515AE",
            x"1EFD84CE6CAA7801F5C68643A479AB28AFE72EE96FCE6399508FCFB6B7C5B424",
            x"2C784F3583ABB402E4A8C9E53EB628EDA7DAE44F07B5956759D7B70083AC067E",
            x"62B4F6C4452906065FAD3EDDDC816D403B825EF68B04751A46930281C52209BD",
            x"1687602EEDEF8909CF21DC088BC301605147CC60D88EA5A3E8FC86C2ADF71E19",
            x"B0CA106440C75F9EB6F28A1DD9A48310DB6BB29105D4BC35CD7BC826A0E2AD27",
            x"093B389EE12A4F6C806EDB28863FC4B900090EFB8C979A44B131BC78B156A1FB",
            x"9FD0D5EC53EBF603C08400EDC95FAF97801F947153F363EF8BCA1AB58B50B2F0",
            x"EF9914C2DDC9E105A1CE0140BF4F2773402F76AB5DEC15C759BB228458598E69",
            x"C767B72608BED38C32B503619E76FA2C606620A848C234AA4610F6CEC4C6558E",
            x"2A1B02F91D9C1D524E8584126DA07362909971ACFD2747ABE93960342F29D454",
            x"6B208677A86A295FF4CC4E3F8030AC16F9E72A2379FA6B29CFD7104666EE96D6",
            x"88F1C9A32C8B6F4FE732F55F4049A23076DAEB7436F388EEB792B8E99844F011",
            x"5D6ABE34E3D80677DACE654E60FE3748A0024826406D5D44837E954E64EF683A",
            x"C90A9D47558409A382359D75917D427DB007FC79E081496FC43CF5759F460C53",
            x"BF9AE96A544E1E35474469247B3967B8080BFAB6D1C37F07AE5B65246E6912DD",
            x"1F624F0BD6F52D456A6E8FFEB0D71B141C19F2801AA43E8B25C01DFE858FBE08",
            x"2E17F6999065E16D0B84D7FC8912A0B62A26EEC022BE5CD8FCA028FCCC571D1C",
            x"6533E0E6789CD301994F13FBDFBEB1816B784420769DCB057BB06D7B32D2A9AA",
            x"9DCDD159B5EB1C826776BDF18F1C8A430834EE70A0E8B88D31088130CE1EAE2B",
            x"68B09B4604C8ABC79A2098EA56ABDBE49C4745A9B14D95D1CB9DC3C9352CA569",
            x"0D89E0690F3DA9AB6371E54BD0A981DFEAEA6C2E0B70749AB968A5BFC5E3BD0F",
            x"905ED08F96D82E28142ADD7999AE428FCA4B82651828A7E2970DBC1FACD51996",
            x"F8CC19D77004656C366A09366625E6D7BBF9479DA46DBBD6F2901A2F2315A670",
            x"75322692280E9D02418B1FC1997CD81311F76B683E8011906EF82366F4B439A9",
            x"25CF78FF6C14E987E258AFA2673B043CBAE2080C5CC03A78847474186786562F",
            x"FCB6357E02374E4BD7C5A7379AD08E5B92571C12CB2053B5CEA6A6249B49D166",
            x"7B81453D074275F993AC3AC36219D5C17FD2AA3E38F0DD04B4B8B97FE07E9B18",
            x"B1436DD98A67A4F67D225224172694A33F9EAB5D5569098F8795973FD0BCE0A4",
            x"8B6400865B9B3F61B9F7DF7E32F8F7B4DF6CA849550F9E574B7472DF999B51BF",
            x"581E01C9C160DE1216E38E3D4E7563070E03ACFF55976DD27826AE0F66605A1F",
            x"442D02BEA3110D3F3055555975A5148A9505237E5472009FB478A5161990C32E",
            x"EE61869CB4BB91DEC8D55547243DB7DAF58DF43DD6AF01EF06B5BDB1267924E5",
            x"C59248EB87917A8C3D15556AFE5803826450E65890A682C68884180BF9B7FF5C",
            x"2C7FFD494B7B32D259B5550A7DC405479ED959C5F9B8C628DDCE2419F603FE4B",
            x"E2BFF97F7830CE1FC605559BB8AE0D6B6C0746ACF615296D08B57E26E105FDF8",
            x"569FF73E3449352FA90D546115A51108020A68A36135EF019D853D78538CF8F5",
            x"50EFE2DD46FFC5E72F915693B43DBB9C071B8DB413C4C682684DD934DD537565",
            x"5947D609687FACDAE77B50FD0658116A0AA150063DAF28C78CF087C7095C251D",
            x"476B911F0CBF23025A30597989C43B0B1AB358095826ED2B5369CBAA9F4A7DA9",
            x"6A097BAE939EF487C348C7365EAE5098A28C441F447841E85C0EB92AEE7BB82F",
            x"0B1F3124FD6C67CBA47D2AC1CCA5D9E5B6D2EE2E6EB4E2CCCA1497EA45B11466",
            x"18AECBFF79029BB93EB9EA22B3BC86DC001E4565848756333B37F3CBEC0BB699",
            x"A5A439FE3786E117DC96CB768D1BC80A002DED1C4FCA514CD0C3EDB9C21900E7",
            x"3C3E56FD434853B38BF03820D1A1BC1B0060C1AAF7BBDB731925C016A727815B",
            x"DA5DD079647CDD0D59E854711A321A208091222A6311802CA7FCA030BAFB4340",
            x"03C898B71EBB099146CCD6ABA34F2371C1FBF76B94BA4063BBFBB04992706461",
            x"85BDE582AC909E7B683310A93476F42AA2F1E2097793E09511F108FE7FA89E93",
            x"4C18DC46A3F9EDB00C4CB9AFC6A0666AB66AD71F237DD1F5BAEB9D7DBF2DECFD",
            x"72250AE8B5F6C00812F39627A8B0998A818A12AEF4389AE4124969381EE0C379",
            x"2F7D9A4D84E0201C3E6D717B2D89E65AC25B3EA46655E25E3FFF0FD42C512437",
            x"E63863F04F50702A5D812B30E05ED9C227C0DCBE99D4D7CD5FFE979662DBFE42",
            x"595495E8F658A86BC843E8C950CC06A77BA10B9CE69713B14FFCF3719601FDE6",
            x"C757F4CD61C5AC89BCE5CD3F593208BA3133996B58F2BD0B77FB6C2A7102F8D9",
            x"AA53E73112AC23DE1B5CB1DE47CF1D934BCD6708456E999823F0026BAB867506",
            x"ABDDDACBBEA2758D204B8A8DEBB6A87C79B11A9CED04E66475E807892949A588",
            x"A98882391CB7A451F0F95AD0C900ACBAB60BA2EB418F599EA4CC0B5FEF7E3C5D",
            x"2E5DC757AB833EDAE97742193F81A392811936486256466CBF32184FC63D5AC8",
            x"65C8AA532944DC024F226727DF42357EC3A7C1FC97D1E9839ECF24F7A959423C",
            x"9CBDABDCEF6F0A07F6F79AFB8E67453C253BA2FBF39ACE456C36FF632F47675A",
            x"EB98298B46069B0BE0636271559A6DDA7DD13671ED6235ED02407E14E66A1A42",
            x"49646E586908E099D09417AB54638083B89BC1AAC11744C187E0BD37598B23E6",
            x"FF1E85C48F9D51E699F63328569541C515E1A22A23B26F224BD199C24658F5D9",
            x"FEACCCAFD7695AD8E6E14CECD0F562ADB4D2376B750F86F7F99A66A7E9C56486",
            x"7CA333A7920F420558537343196516A0071F420825974863F66398BBCEAD1FC8",
            x"BBB4CD3B7F16670D44DC2C64A71DB0B00AAE671C7C727C95E1956591B4A1AFBC",
            x"910731D03EB19A916F0A629FBAA809881AA59AAABAAFBBF4D2751C7A07B2271B",
            x"7B8ACA985C8A62FB069B96EF12AC1E5C22BC62AA92A711E71FA5AAB30B0F7AA1",
            x"315A3AE4CBDB967088E17046BEA22DCA769A96AAFEBABADAAF3C2A8C989632B3",
            x"CB43525F398171A9DD5328E89CB760BBA0E2F0AA7C929202A6DA6AD3E5F14E8C",
            x"38645FCED6432A2E895CED4DEB821191315669ABBBFEFF06B8038A1DDCEB74D3",
            x"D49ECFB411E4EB64DF4B4170C9473A7BCB518E2911FC7E8894055B288B48271C",
            x"17EC37063ADF481F0E7863293F6AD3B1B85A556FBAFABCDDF60D40EDD87C7AAB",
            x"B3C24289520E7C2E95B494EFDE0A1D0A14C3D50712729B08E111614084BAB2A8",
            x"8DA7E6DF5F15BA64F407F7478D1B299B3725958ABFAEE09D53BB1361CF928EAD",
            x"503BD80E4EB4139F660BE26B51A0EE60C2FC745A9F2451E95D10BC12B77ED4A0",
            x"D8518415F4863D6E1919D7885A314591267AA6C2EEFEDACF49B99A3E823C17B0",
            x"04DA4E34E7C9590527A6935CC34B6C7BF9B2B826447C02367E16635CC75A3309",
            x"8F03F5475BBF478DFB38FC4B247802B1F60E9479EEBA0741BD31944B2A434C9F",
            x"5685E56A411E6B50F0D57AF8FEB4068AE114F6B6C4930A6219CA76F8EBE473EF",
            x"50CCDD0BE3AD8859691532757C8608DA53B760802FFC9B9726BBA07549DEADC6",
            x"D9330999D5205CC70FB5CFA53BC91D03DD0211C067FBE172F89130A57E8CA0A9",
            x"87CC9E6695F0CB2A9704B73DD1BFA98589873AA09BF1D32E75FBC9BD3CD3B1AE",
            x"CBB3ED98F4E938EAF28F82D89A1F2E4C5E4AD2B1E1EA9CE5A4F1BE19DB1D0A24"
        );


    type casr90150h_vectors_t is array (0 to n_gen_rand-1) of std_logic_vector(511 downto 0);
    constant casr90150h_vectors : casr90150h_vectors_t := (
            x"ECCE6F82DF3C15F90368B1912179107C28EC63F150681C1CDDF8A19F05B54D682E9F41C01F344725FE31A6F40414DA6BC1FCF9D36AF8D942701992609FA010D9",
            x"C3B5854416EA35CE840D2AEAF33FA8824D8E944A18AC3E3BC1B512E48D117C0C626E63E023E6E8FCD54B9C260E2783EA63C37F8F68CD8767D8267FD165303946",
            x"26844D6E20EB45B84E11C2827CD50DC5F4D8F2FB250269426305AEDFD8AB2612D5A5B690743865631572FE7B1759C5A9F4A534596DB8C83BD47BFBDB3DC8562A",
            x"7A4EF12F71E96D2CF53A6647AB9595ADC3CD6ED1FC85EE25D58C8485DDA8FF3CC19CB2E8E274BD16B52CC9FAA056280F079CC6DE60ADBC71C6B3B1C2F0B49749",
            x"31F46BCC3A6E08CFD5D3F9AE29F46109A57D009B3B4CA17D55534F4CD12D61DBE3EB3C0D97C7B1A2A5EFBEB8B0C34C118A732A13F108BA8AE80F0AE4C987753F",
            x"CB668BBA4BA5153A041D1EA96E66F29719758161D3739268141E367B4AE513031668E214F66A2A349CC8A89D99A6763BDB9DE12E9B95305A2C149A1BB64B60FC",
            x"3B18DB39F19CB4EB0E29A426059A1EE1A76042335F1F6FCC362F71BA3019AF86A7ADF523A5EB4157E3350DE0769B85724071D2EAF3E5E8C34237E323A3F1511B",
            x"D3A502FEFAFB8761956E9E7D0CE938731E50E76D0DBC627241645A99583628CA3C8054F5B9296341F4C09490F273C94DA09B9C401F7C6DA4274194F797EA1AA2",
            x"1EBD84566AC04933E50465E493C7E49FA9995F2091AAF7FDA25E926F1C5565B94F40C7309ECE3662C72163F93D9F3F3591F862E03C02A09E5B627325F1C32094",
            x"2E184ED382A0F6FC7D8EFC1BED29BBF40EEF4BD17B881629B78E6F8CB28119973161A9D960F563942AF235BFC8FCFAE1FBCC94506A06116D9115ECF84AA5F1F6",
            x"6724F61F4611624688D49238C1E620D6108A781A72DC256F8257E7DB9CC3BFF0DA3287D751843766426D7015FDCBD23310BBF6C8E9093B206AB48734F0BD2B83",
            x"19FF6324692A15EC5D977F4D225B51033953B423EC9A5844C7913B0B73650069D16E48C61BCE601BE78C1834A83B1F6FB9A8E2352F97F2D0EA07CEC3C990EA46",
            x"277E16DE87CB35EED8F2563CF7CA0A87F71D0254037194AFEA7BE0927F59808E4A25F56D2875B03BFB5E3447AC62AA60B7055550C5E34C992B09F067367989AB",
            x"F93D3206CB39C5E895EF914773311AC8C6A587D6071A632403F3317DE5164157B95C5445E4C5284BD84372A922B40BF1238C54496C747367C99EA8DCE3BFDF0A",
            x"76D9CD0A30E7ADE56447FB2F3CCBB2352C384E1109B1F5FE04AEFB309CA5E251864AC6A81BECC4F38CE71EA7F436198AD45AD6F662968E3BFFEEAD4FF7164998",
            x"A286B19159FA29F83EEB18EBCBB33F74C65CF13A9FBA912F0FA680C9F3B8D5DACFFAAAAC28232F7F5B5DB8B9B6732658D6DA1277F46057718E46A53140B1BF64",
            x"B4488A7B5E4367CC6CC8AD80B98EEB172D876AF26CA0EAE59E3A41B6BE050100F05200A66455CC244845A59E139EDD85D01B3DB496B0D00A55EAB9CB618B997F",
            x"06FDD99A55E518BEA3BD08C186DE29A1C4CE0ACFC3112A9DE551A28287098281B8DF01BDDA95BA7EF4E998672FFE8C495839D113E239981B854896FA3250E65D",
            x"8AF88669C47CADA0159995E348874F13ABF91AB667ABCA791C1A9644C99E4442858E830C4A7539A64747F4D8E54E56BE046F9AAEB56EE4214C7DF4316DD99F89",
            x"58F5CBA6AE8BA91024E6F4157D4833AE093FA221D88BFBE6A22061EF7779EAE449D44796B3C4FE3BEA6C534D1D77D4BB0EAE68AAB52CFE5332B8A24B288FE85E",
            x"C5E4BB1AAC5826A85FD8862029747C0F1FD33753455B801A3770F24C7166C0DEBF16E8640C6F574BE38ECC39B91113B3948D85A0B5CBDFDCFE15B7BAC5DE0C8F",
            x"AD5F92A8AAD47A84DF0549706F26CE1DAB5CC75D2C53403143699FFAFA5C218E09B0E4DA1EE75073F55AB65E07ABBD2EF7D94D31B4310D0B0D340710AC8517D5",
            x"204F7C85A286B8CB9E8D377886FA713108072F48E2CE205A254EFF78299E73D71FA9FF5320BB58BFC5483587098BBDC2829E78DB367B919890C60EB90BCCB4D4",
            x"70F63BCC36489D30FC51E26DC8F9DAFA9C0EE37D94B750917C368E3C6779BE10B88E450CF1314D85AD7470489EDBBCE446F5BD1BF389FAE5E9AB109793BB0356",
            x"A9E153BA51FDE0F9CADA37CDBDFED248EE185519F730096A72425552D96603390555EC97AAEA784C092298B5FE93BF3AA85510BA9FD650FCAFAAB9F5FF198713",
            x"2F535F39CA49D14F3A83637D08764FF5612CD0A721F81E49EFA5855C5E5D07D788546BE7A2AB9CFA17F47584AE6FBAF00CC4B988FD01D9DB86A896A054AFCDBF",
            x"E55C4CFEB3FF9A7BE24474649CA3B2D433EF191BF34439BF0E3CCD42979D8C11DCD6A29FB608636933E2904FA7A5B208132F9F5509820601482DF4B0D7AE753C",
            x"5C4AF3569D4E698877EEC6DBFB373E066D0AA6A02F6E678D9D5BF164E07C5E3A5F9014FB851CB607EDD468BD399CAF1C3DCE65409EC70B033C60A389912DE0FB",
            x"4AFA6E52F17587549344E8D8E0C0E90BA592BC106527FED1E0031B1F10EED35198F82721C8ABA309E892AD91C6FB02AE79BD9C61FEAA9A84EA91B55EFBE91112",
            x"F8F387DC7B1549436C6FA5DD51A12E9218FE9E38DCD988CB1006B0A4A9000F5AF5D459F275081696E5FC047AEAC28683D72162938E02604F2A7A010ADBC6BABD",
            x"F5ED4982A8A4766522879C544AB3C0ED25B0E975CB965DFBB80A393FA6801940B116DFBFE09C32E27CF60AF808A44CC653D214EE5707B0F6CBB103988BA810B8",
            x"65417E44A51EA3B8D64BE282FA0FE168D8894E057AE39D229C1967D53AC03E611AB0940B116A6C5593671A3C1D1EF76F9C8F374B808BA9C0788B8565532439B5",
            x"1C633FEFBDBCB62D81F93646631DB2250557710C70F77CF462277B15C8604393B0296618BA6BAAC47C1DB35239BEC660EBDFC17241518E20C55B49595EFE5725",
            x"AA94DDED00AB834DC277E1AD94A03F5C89162A92E9D04FB6D77840B4F4D0E6FF984F3B351BE8002E9225BC1D46AEADF1A896A23DA34AD7516C423F07467595DD",
            x"287708E98108477D27A332AD67306B53DFB56A7E8F08B292D374A10737495EFDF4F6EBD1A82C006EFF79AE212A06048B8DE0B5451672905B62E55A8C6BA5F1C8",
            x"6CA29D66439CE904DBB4EE2C1AC8E94E8B810B9C559DBE6CDD671388D13F52F833C0E2CAA442008E563F8173E90B0BDAD1F18468A39E78C076DD02D6A33D2BFC",
            x"8336E93BE5FB468B9187AD6E32B52E7ED9C398EA95F829C3C058ADD54ACA4CF45E21F47A3AA701DFD150C36F8F9A99C0DBDB4E8597F595A0D089865616D0EA9A",
            x"C7C04FFBDC416AD0EACB89495E05C186066565EA75444F6660850015307BFFE69B5256E35A1B82959B59A44D55F066E1C0997EC96154F491495E4D97321988E0",
            x"2820F5DB92E20009EAB9D7365D0CE34B0DD9196BE46EB35BD1CD8035D8E1E05A735FC2140B2044E4684F9AB90458BC3361FE36367347C77B3E4FB474ED2FDD31",
            x"EC71648B6EF700176A1652D5D99B3573944FA6281EA6BD125BF0C044DD12D0C1FF4F252211D0EF5EA4F8F29F8ED53E6F73C54357DE6B2810EDF502E3E9EE4CEB",
            x"C2AB1FD20CD380272B319EC196EAF01E72BB3D4C2E1AACAD88A9E0EF50AE09A22976DCF73B596C569F7DDEE55685F9E14CAC6744DFA0CC392165861766CDB72B",
            x"A428AD9D1B8C405FC8CAE4E360C018378E18DC7267308721D5AE31CC09A117B56E009336D9062AC2E635181D024C56B2338A996B5D91B277D21C4D343A3985CB",
            x"3E6DA061B9D2E0D23DBABF9511A03470512D0E8FD9F9CFF355277A3A1733A48543016FD4CE8940247940B42185F2D4AD6C52EE0318EAAD83CF2AB5C2795FC9FB",
            x"DF8030B20E0E510F689237E0AAB07298DBED90564746F23F14F8435921DD3B4D27832CC3F85E607E9F6132724C5C938462CE4F07B5E200C5F7E880E59F467F92",
            x"0CC049AD1D15DA9B2D7F6311AA08DEFD010C78D1A96A1F4DB734A44FF3DDCB71FCC4CB653C8DB0A6E612FFEDB2DB7D4AF63DFD8C347701AC924DC118E469F87C",
            x"13A0FE09B1A588F9C13E74AB2B155840839EB59BAE293B3183C71EFDBEDCB32A2FAFB359D75129BA793CCB881C921D388161F15E76928283EFF0E3A5FE8734DA",
            x"3EB17F161A9D554F23DDC721E8B514E1C5E081E0A74FE1DBC4E8BCF0065F9FE96087BF16571AC6099FD7B9543B6D2DF54233EA53D26E4445A669153856CBC341",
            x"DE0B3CB33A78547BD5086AF3CD05A373A811C3713975B3526F0D2BE80B9B704F514BA5A597A22B166794A7164221C480277CC1CECDADEEEC198FB1D4D2306723",
            x"8F18DBAECB84D688059CE2BCB18C151E0C3AA50AD6143D0DCF91C944127038F40A799D38F69742A3BB731EB3A5522BC05B0323BA708866E237D50AD39D48DDD7",
            x"55A5030E31CF12D40CEBB6079ADA20B7165AB89AD3266C917E7A7F6E2DF84DE61996F0C5A47364B7382FB88F3D4D49E08185F609D954BAF772159A5FE175CDD1",
            x"55BD869F5A37BC0213C9A10E728951B1B58A9562DFDBE76A75F1CE0F69A4FD5B37F0D968BACD3F90FC68A5DCC9717EB1434DE317D74730C25F346389732575DB",
            x"55984AE45B7212072D3E9399BE570B3B20D2F036CC13BF49E5AA751C473B6442D4499E4D1AF0F569528518C37F1B18AA2579D7A4C06AE9A79FC6D55F0EFC61C2",
            x"D5E4F87ED81F3D0FC1DC7DFF0DD099EBD1DE6860F22F2B3F1D29D5A2A9C01AE4C2FEF7B5AA8945075EC8B5666CB2A5895C0F903B60A2EE9B7E2A51089E72D3E5",
            x"955F74961C3FD09A220AD0239019F7E29A418CB1AD44C9CDA0EE44B4A7E038DFE4DCD010A25E6D884435315BC33C185E0A1E784B7116E6604D699B9D67AEDEBC",
            x"F44E27F3326E99FB571AD874682E96F4E3A2572BA06F7F71B107AF07B8904D8D1B8B8829378DA854EE40FB0BE6EA248B1B35BCF35BA0FBB0B00E616D392CCABB",
            x"E6F579CEDFA4EFC942A2CCF28C6EE45775B7D7C8B0A44B7B8A8986890DE8FDD1B2D9D46FC6D104C76DE1C0939AE95BDBA1F5137F1391D3A9B817D345FFEBF8B3",
            x"DAE536BE179F4CB66636FBBED28E3AC10087963D091EB962D2DEC857998D651A9C8606C36CDA8F2828D321FF70EF41C293D4BF21AFEA1F8E2431DC2855C035AF",
            x"80DDC2B723FF7BB5B94099800E5F6222814F75789EBEA654DE4EFCD17F5518A07F490A644FC2DCE4451FD2B479E462E47C8795F305632DD55E4ACE6CD4A04105",
            x"4188A4A0F54F3A31A7616EC015C47754C33A20156E2E9D87C5B68B9B6501BD30E97F91DABA66035EEDA00E86E67EB63ADBCA75FF8D34C0151DF871C797B0A28C",
            x"E3DDBF917577D97B9A136CE0242ED74724DB70344746FDC86D0259EA5C8204C98E1FEBD21BF90656683010CA1B8E2570C0B3A5E051F7A035B974EAEDF10934D2",
            x"56081D7B35128E08F33C6B907E6E4769DBC82866A96A0D7CC885964193C70BBED32F62CF28168BC3A448297133D75949E1BC3DD08A53906426270A044B96C35C",
            x"D31C291AD5AEDF15DCDAE1E8AD8FAF2781746CB82E29146BF5CCE1E26EEE929ECFC63472E430D3A71EF44F6BDF00473F33225189D9CDF8BE59789B0AF370E70A",
            x"1FAA6FA8048405A11B82B205A0DD03D843628734674FA2CA25F3B255CE00EC6EF02976FE9A691F38A462F243DC80EEF9EDD7DB57D638553D9635E098CE299D98",
            x"2CAB85040F4E0D12B1C62F093181849CE456CFE6D97516F97DAFBFD4FF014E86B84F12286BEEA4CD9E94DFA7DB41E01721828B44C36CD5F8614491E5BF67ED64",
            x"63294D8E1E7518AE3A294E96DAC24BF37A943278C615A4A67125AF1725837A4A04F6AD6CC0249F3864F39B39D2627035D346D36B662B9454F26FFA98B41A047E",
            x"97EF705F3594AD89636F3C6412A5B8DF12724F95EB241B3BEAFC86B0FD4429F90BC00847E05FE4CCBF6EF0DECDB588615D681F037B41F6D71F85B2E5262B0ADF",
            x"704628C4D4E7A9563406F2DA2E3C2515BFEFF2F50BDE31C2023B4809202A67779A2014AF108EFF3BB60AD94670B4DCF20824258742624292BECC0E19DB61984D",
            x"28E96D2F07FA264576088EDB655258A53B0BEEC49A1F7B6507523C17F06B9D21F15027A2B95454CB2110972BF9378F0D1C5E7D4D25B7E47EACB211260A13E4B1",
            x"EDCF01CC8B437BE8111D5CD91D5D959CF091C0AF613C415C8B1D6A31B8C974F23A5858361E16D732D3B966E3A7F1D294AAD5B07CDCB37E9C830D3BFF113C1BAB",
            x"C13682BBD0653AE42BA903DEB9406173497AA10752EAA21B51A96B4A0D7F33ED41C4DC55213010DC1D1E3C17395A1EF30A0508A75B3C1E6BC591D1B8BBD2220B",
            x"A2C0C4BB88BCD87A49AF85508760F21F7F7AB28B1CE897331B2F6871186ADE41232F9281F2E8391221A36E30C751280F9B0C95BD12E22FA9EDFADA153B9F751B",
            x"34A12FBB552B0C8BFEA7CD09CA111F351A7A8E59ABEDE7DFA9E46CABBCCA13E3F7C7ECC22EAC7FAD52372149684BCC10E19BF504ACF7458EA1704331FB6760A3",
            x"C733E53A45C99BD04C3B7997BB3BBBF4A3FAD1C7AA60BE5CA79EE323037B2E57342B6B67680295295F45D3374CFB3639B378E48B83D26CD49228A4CA5A1B5196",
            x"29CDDDF9EC3F6A88F2505EE600DB20D7953A1B2AA9B1A99B3A6EB4F68760EBD0D248235E4406F5E746690CC033C2E577AD0D5FD2470FA397EF6DBB79C9291B72",
            x"6F3088DECA6F00D5DFD8849D018AD10071DB21CA2FBA0FF3DBC637E2C9514219CDFC5719AA0844D8698697605F24F9448098448DA89F97F3A700107637E6A34D",
            x"05C9DD0633A781011F054F7482D04A808A48F33B64A1123E48EB7354760B6526755AC1B6A31CEF1CA64E66509CDFD72B41FCEFDD0D77F14D1B8038E761D83731",
            x"8D3E898B5D9A4282BE8D3E73C698BAC1DBB56DF15F13AF4FB50A5C56F31818FBF042A31435AB6CB399FBBD99FB9D16CB23C34C9491134B71B0C0551C328C45EB",
            x"50DCDE5250F3E4C62C51F5FCA86DA2238181054A0DAF033484999AD23FB43DF338E617A241892B9F6EFAAC6EA3F9B47BD4A57BE3EBAC7A0A39A091AE6CDAA9AB",
            x"598B0FDDC9DCDF2D42DA0427AC88175642C3887B118485D74FE6F29D4412456EC5F92037A3DEC3742C7806CEB746A2D2579C3AD6AB8A911B67B1FA23AB0A2F0A",
            x"C7D89580B61B05CC66830E7E23542743E6E55C91BBCFC9413E9A9E612E2FE806E957D057B44C26364ABC0C7E906A165D927258068BD27BA07A8AB37782936199",
            x"A805F44191318DBEB8449DE174565F66FC994F7B9235FE22D4E07D93EF63C40A8E53088782B25B53F29616F6E8A9358DFF9FCC0EDB0F9390C2588C65C4FD5366",
            x"AC0CE6E26BFB592024EF601236D39B3A5F6F7310FD748974D710C8FF8D55AA1853DC95CFC62FCA4FCEF724220D0FE0551E76BA1A529FFFF967C5D6D82F701F7A",
            x"A2135A7581414ED05FC6702F509F71E9CA4A2DB9B817DE77D3B9FDF5580021248E0B65F36D46B1FDBC65DA7511957090AD9099398C775D577A2CD4444C282950",
            x"B53C418443627E08DF29C86B49645BE7BBB365B79421D9F05C1608651C0072FF53183DBC4C28AAE0329913E5AAE509F90169EECF52924952436352AAFA646E19",
            x"04DAE24EE437B7159EEE74C17F1E90F8318C19A2F652D73882331C9DB200BCFC0FA4610EBE4D80506EEEAD9C28FD9E968227CE390C6FFF5FA5161EA8D99EC326",
            x"0F8255FE5E7201A1FCC5C7E22EA6E94C6ADE2796A3CC47C5474EBB601D0187FA109EB29011B140C8AC4A04626DC8E8F6475ABF4E92AF5C4F1CB328AD8E64E7DB",
            x"94C7D4D7D59F03134BAC6B17643A2E7AAAC17EF03632AE6C2B36201030824C71296C3CE83BAA61358AF10AD5C03DED07AB5A957AEC0E4AF6BB0EEDA4DF9F9CC2",
            x"F7AB971184FF87AD79A2E0A71E5941888AE338C8437C81C261C3503859C7FEABEE22630C588BB3D4526A9A54E068658C895AF428221DF8C0A196043B8566EF64",
            x"60A970BA4FCE480C06B6B13FBDCF2355DA94D5BCA70BC365D3E6085C9FEFE22B0357B7968D582F86DF80739710ACB8575E5A6664553055A193F30A53CD18817F",
            x"112F29B9FF35F41E08002BC2083CD545827311BB399BE55D5C9B1CC3F483D56A8753B0645C044D4A07409D70A90334950DDB9B9A85F8D4926C6E9B9F39AD425C",
            x"3AE6EE3EE6F5E6311C0041671C53406D47ECBBB1D7F3B81803E2BBA7B7C580084D5DB8DA860EF9710A617D69AF86E3F091986A78CC4D977FE286E168FE28258A",
            x"50D8477658D5DB7ABA00A35FBADE20A86F0F90AB505F2434049421B910E8401CB448AD524D145F3B93920D4625CAF5897B7C81AD72F8F01FB64A134DD7647959",
            x"5984E803DD858B0A2301141202875184A29B790918DCDA560FF6529FA90CE02B12FD080FBCB6C4CB7D7D152B7C38C05E5103C32C5CCDC82F31F93C34101EF607",
            x"47CF4C0790CD53935483B62F06480B4F9668369EA59B53831EA38E652697506AACD9941397202F321134A1E26A65A08B9A84A7EE9BB83C46FB77DE423824A708",
            x"E836720969B05E6D4745A16B89F4197C75C4446C3DF20CC7A4B7D59DFAE648882786E62DF7D04CDD3BC31295C9BC91DAE2CFB8CAF3AC7AE80121C9A57C7F3D9C",
            x"4C41AD1706B8C7AC6A6C93405E663602806AEAA2595D17E8BF8144E0A81DF55C7CC8FB642658FB11F9A7AEF4FEAB7AC0B63E1D301F8A90EC02F2FE3912B7DD6B",
            x"72E221B08825280EAB837C20DD9B7504C0C24A178659A60D16432FD1A43CF04AEFBDCB5A7D855AAADE3C80272E0A1261216520D83DD279E206EC3957BC824C6A",
            x"ACD77229D45CE41809C4527118EA508F21E7FB32CBD61D10B1A6C71A3E4F78F880B83313F5CC48A005574078E7193FF2D23CF11C680F967708C25715B3C7B6E9",
            x"23922D4686DB5E3C1E2E9FFAB5C189DDD21FF1EEFA033CA90B3AEAA947B22DF541347FAD2172F5B00D5560FD18B7FB8CDF636AB6EC1FF3829DA596B0AFAA862E",
            x"76FF616AC89147663D64672A94225F919F23EB64B106EF2E91D0AA27281F6D6522E68425F24E441819503131B5315157CF35009622374FC6F9BC74890D224F47"
        );


end package casr_test_vectors_pkg;

package body casr_test_vectors_pkg is

end package body casr_test_vectors_pkg;